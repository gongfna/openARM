//
// cortex-m0-nvic.v
//
// the nested vectored interrupt controller for the cortex-m0 cpu complex
//
// Danny Gale
// 9/15/2016
//

module cortex_m0_nvic (
   input clk,
   input reset,

   input [N_EXT_INT-1:0] ext_int,
   input nmi

   // needs a bus interface
);


endmodule;
